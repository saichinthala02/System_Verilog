mailbox mbox=new(); 
class eth_pkt;
	rand bit[55:0]preamble;
	rand bit[15:0]sof;
	rand bit[41:0]sa;
	rand bit[41:0]da;
	rand bit[15:0]len;
	rand byte payload[$];

	function void print(string str="Eth-Pkt");
		$display("----------> %0s <-------------",str);
		$display("preamble:- %b",preamble);
		$display("sof:- %b",sof);
		$display("sa:- %b",sa);
		$display("da:- %b",da);
		$display("len:- %b",len);
		$display("payload:- %p",payload);
	endfunction

	constraint l_c{
		len inside {[10:15]};
		payload.size()==len;
	}
endclass

class eth_gen;
	eth_pkt pkt;

	task run();
		repeat(10)begin
		pkt=new();
			pkt.randomize();
			pkt.print("Eth_gen");
			mbox.put(pkt);
		end
	endtask
endclass

class eth_bfm;
	eth_pkt pkt;
	task run();
		forever begin
			mbox.get(pkt);
			pkt.print("eth_bfm");
		end
	endtask
endclass

class eth_env;
	eth_gen gen;
	eth_bfm bfm;

	task run();
		gen = new();
		bfm = new();

		fork
			gen.run();
			bfm.run();
		join
	endtask
endclass

module top;
	eth_env env;
	initial begin
		env=new();
		env.run();
	end
endmodule

/*
# ----------> Eth_gen <-------------
# preamble:- 10010010101001111101100011000011111100001001101001010111
# sof:- 0010011111011101
# sa:- 111111010101101010111101111100110101001101
# da:- 010010001111100011000001101001011011001001
# len:- 0000000000001100
# payload:- '{71, 55, 66, 124, -71, 106, -67, 15, 98, -80, -80, 2}
# ----------> Eth_gen <-------------
# preamble:- 11001110101110010011111101011001101000011001101110111110
# sof:- 1111011000100110
# sa:- 111011111111101011100000010111000011101100
# da:- 100011010000011011000111000101111100011000
# len:- 0000000000001110
# payload:- '{-108, -72, -56, 90, -96, 55, -71, 122, 54, 73, 95, -126, -86, -22}
# ----------> Eth_gen <-------------
# preamble:- 11100010001010000000000001010101111001000110000000110101
# sof:- 1111100110110110
# sa:- 111100001011000100110110000000111010100110
# da:- 100110001111000111011110101100011100010010
# len:- 0000000000001101
# payload:- '{70, 18, 107, 78, 120, 50, -90, 72, -83, -65, -87, -122, -71}
# ----------> Eth_gen <-------------
# preamble:- 01110101111010101010010011011011110111011110000101000011
# sof:- 0110001001011010
# sa:- 110101100111011110001111001100110110101100
# da:- 111110111100011101001110101000111111110111
# len:- 0000000000001010
# payload:- '{74, 69, -115, 102, -21, 23, -123, -127, 63, -43}
# ----------> Eth_gen <-------------
# preamble:- 10001100111101010100011001000010110100000010000100010100
# sof:- 1110000000100010
# sa:- 000101011011010001000010101001110010000001
# da:- 010010001000101111001011100011000000110111
# len:- 0000000000001101
# payload:- '{12, 62, -111, -16, 41, -113, -41, -77, 11, 48, -51, 28, 115}
# ----------> Eth_gen <-------------
# preamble:- 11000111001000010001010010110000100100001101101100100010
# sof:- 0101000110100101
# sa:- 111011000000110010111011010001010011110101
# da:- 111110000100111100001110011100010101100000
# len:- 0000000000001111
# payload:- '{-35, -6, -31, -23, -66, -31, 53, 81, 23, -30, -49, 100, -81, 20, 111}
# ----------> Eth_gen <-------------
# preamble:- 11110110111010101111011101011100000011100101100100101011
# sof:- 1011100010001000
# sa:- 101100011100111100100111101010001100011000
# da:- 111110110101010110011100100001011111011010
# len:- 0000000000001100
# payload:- '{-18, 117, 4, -33, -114, 58, -114, -11, -19, -88, 44, 88}
# ----------> Eth_gen <-------------
# preamble:- 11110001101000101000000111011011000111111001011101011001
# sof:- 0100111110000000
# sa:- 111101011011110101011100011101011110100110
# da:- 010000001011111000100000001111100000001000
# len:- 0000000000001010
# payload:- '{-117, -72, 32, -54, 125, 28, -65, 73, 63, 105}
# ----------> Eth_gen <-------------
# preamble:- 00011010100010101010000001011011111011011010101101111111
# sof:- 1010011100000110
# sa:- 101100000100000001101100110101111001010000
# da:- 110011100111100101010010111101100011001111
# len:- 0000000000001110
# payload:- '{61, -22, -100, -98, -37, 97, 94, -49, 9, -24, -64, 35, -95, -38}
# ----------> Eth_gen <-------------
# preamble:- 10001010110011100110101000111010110010001100000010110100
# sof:- 1001111000011000
# sa:- 110101010001011110001011111110111000011001
# da:- 101100001110100100101010100101100011100111
# len:- 0000000000001011
# payload:- '{-49, 87, -27, -49, -11, -35, 60, -4, 95, 61, -55}
# ----------> eth_bfm <-------------
# preamble:- 10010010101001111101100011000011111100001001101001010111
# sof:- 0010011111011101
# sa:- 111111010101101010111101111100110101001101
# da:- 010010001111100011000001101001011011001001
# len:- 0000000000001100
# payload:- '{71, 55, 66, 124, -71, 106, -67, 15, 98, -80, -80, 2}
# ----------> eth_bfm <-------------
# preamble:- 11001110101110010011111101011001101000011001101110111110
# sof:- 1111011000100110
# sa:- 111011111111101011100000010111000011101100
# da:- 100011010000011011000111000101111100011000
# len:- 0000000000001110
# payload:- '{-108, -72, -56, 90, -96, 55, -71, 122, 54, 73, 95, -126, -86, -22}
# ----------> eth_bfm <-------------
# preamble:- 11100010001010000000000001010101111001000110000000110101
# sof:- 1111100110110110
# sa:- 111100001011000100110110000000111010100110
# da:- 100110001111000111011110101100011100010010
# len:- 0000000000001101
# payload:- '{70, 18, 107, 78, 120, 50, -90, 72, -83, -65, -87, -122, -71}
# ----------> eth_bfm <-------------
# preamble:- 01110101111010101010010011011011110111011110000101000011
# sof:- 0110001001011010
# sa:- 110101100111011110001111001100110110101100
# da:- 111110111100011101001110101000111111110111
# len:- 0000000000001010
# payload:- '{74, 69, -115, 102, -21, 23, -123, -127, 63, -43}
# ----------> eth_bfm <-------------
# preamble:- 10001100111101010100011001000010110100000010000100010100
# sof:- 1110000000100010
# sa:- 000101011011010001000010101001110010000001
# da:- 010010001000101111001011100011000000110111
# len:- 0000000000001101
# payload:- '{12, 62, -111, -16, 41, -113, -41, -77, 11, 48, -51, 28, 115}
# ----------> eth_bfm <-------------
# preamble:- 11000111001000010001010010110000100100001101101100100010
# sof:- 0101000110100101
# sa:- 111011000000110010111011010001010011110101
# da:- 111110000100111100001110011100010101100000
# len:- 0000000000001111
# payload:- '{-35, -6, -31, -23, -66, -31, 53, 81, 23, -30, -49, 100, -81, 20, 111}
# ----------> eth_bfm <-------------
# preamble:- 11110110111010101111011101011100000011100101100100101011
# sof:- 1011100010001000
# sa:- 101100011100111100100111101010001100011000
# da:- 111110110101010110011100100001011111011010
# len:- 0000000000001100
# payload:- '{-18, 117, 4, -33, -114, 58, -114, -11, -19, -88, 44, 88}
# ----------> eth_bfm <-------------
# preamble:- 11110001101000101000000111011011000111111001011101011001
# sof:- 0100111110000000
# sa:- 111101011011110101011100011101011110100110
# da:- 010000001011111000100000001111100000001000
# len:- 0000000000001010
# payload:- '{-117, -72, 32, -54, 125, 28, -65, 73, 63, 105}
# ----------> eth_bfm <-------------
# preamble:- 00011010100010101010000001011011111011011010101101111111
# sof:- 1010011100000110
# sa:- 101100000100000001101100110101111001010000
# da:- 110011100111100101010010111101100011001111
# len:- 0000000000001110
# payload:- '{61, -22, -100, -98, -37, 97, 94, -49, 9, -24, -64, 35, -95, -38}
# ----------> eth_bfm <-------------
# preamble:- 10001010110011100110101000111010110010001100000010110100
# sof:- 1001111000011000
# sa:- 110101010001011110001011111110111000011001
# da:- 101100001110100100101010100101100011100111
# len:- 0000000000001011
# payload:- '{-49, 87, -27, -49, -11, -35, 60, -4, 95, 61, -55}
*/
